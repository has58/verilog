module new(a, b, a1, a2);
	inout a, b;
	

	assign a= a|b;
	assign a= |b;

endmodule
